///////////////////////////////////////////////////////////////////////////////////
// [Filename]       -
// [Project]        -
// [Author]         -
// [Language]       -
// [Created]        -
// [Description]    -
// [Notes]          -
// [Status]         -
///////////////////////////////////////////////////////////////////////////////////

module rom_cordic #(
    parameter int Width = 16
) (
    input  logic [      3:0] addr_i,
    output logic [Width-1:0] data_o
);

  always_comb begin
    case (addr_i)
      4'd0:    data_o = 16'b0010110100000000;  // 45.00000000 45.00000000
      4'd1:    data_o = 16'b0001101010010001;  // 26.56505118 26.56640625
      4'd2:    data_o = 16'b0000111000001001;  // 14.03624347 14.03515625
      4'd3:    data_o = 16'b0000011100100000;  // 7.12501635  7.12500000
      4'd4:    data_o = 16'b0000001110010100;  // 3.57633437  3.57812500
      4'd5:    data_o = 16'b0000000111001010;  // 1.78991061  1.78906250
      4'd6:    data_o = 16'b0000000011100101;  // 0.89517371  0.89453125
      4'd7:    data_o = 16'b0000000001110011;  // 0.44761417  0.44921875
      4'd8:    data_o = 16'b0000000000111001;  // 0.22381050  0.22265625
      4'd9:    data_o = 16'b0000000000011101;  // 0.11190568  0.11328125
      4'd10:   data_o = 16'b0000000000001110;  // 0.05595289  0.05468750
      4'd11:   data_o = 16'b0000000000000111;  // 0.02797645  0.02734375
      4'd12:   data_o = 16'b0000000000000100;  // 0.01398823  0.01562500
      4'd13:   data_o = 16'b0000000000000010;  // 0.00699411  0.00781250
      4'd14:   data_o = 16'b0000000000000001;  // 0.00349706  0.00390625
      4'd15:   data_o = 16'b0000000000000000;  // 0.00174853  0.00000000
      default: data_o = 'x;
    endcase
  end

endmodule
